��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  A�Z�    PAR      �  )AQO    SUMA2      �  1�Y�    SUMA1      �  a	�    X2'+X4'      �  Y���    X1xorX3      �  � (    CARRY      �  Yi}w    X1+X3      �  Y1w?    X2X4      �  Y� w�     X1X3      �  � q 
     X4      �  � q �      X3      �  � q �      X2      �  I q Z      X1                    ��� 	 CLogicOut�� 	 CTerminal  L�a�              @            <�L�         ��    �� 	 CInverter�  `ha}       	        �          �  `�a�      	       @            T|l�          ��    ��  `hui      	        �            t`�p           ��    ��  `�u�      	        �            t���     !      ��    ��  0E      	        �            DT      #      ��    ��  CXOR�   `5a                          �   p5q                          �  Lhai               �            4\Lt     &      ��    ��  COR�   �5�               �          �   �5�               �          �  L�a�               �            4�L�     +      ��    ��  �(�)               �          �  �(�)              @            ��4     /      ��    ��  CAND�  �(�)      	       @          �  �8�9     
          �          �  0!1               �            �$<     3      ��    1��  ����               �          �  ����              @          �  ����               �            ����     7      ��    )��  P�e�              @          �  P e              @          �  |���              @            d�|     ;      ��    $��  P�e�                          �  P�e�                          �  |���               �            d�|�     ?      ��    )��  �     	          �          �  � !               �          �  1               �            $     C      ��    )��  P�e�                          �  P�e�                          �  |���               �            d||�     G      ��    1��  �P�Q     
          �          �  �`�a               �          �  �X�Y               �            �L�d     K      ��    1��  HH]I                          �  HX]Y                          �  tP�Q     
          �            \Dt\     O      ��    1��  H]                          �  H ]!                          �  t�     	          �            \t$     S      ��    ��  0� 1�                            �  0� 1�               @            $� <�     W      ��    ��  � � � �                            �  � � � �               @            � � � �     Z      ��    ��  CLogicIn�� 	 CLatchKey  � � �       ]   �  � �                             � �     `    ����     \�^�  � � � �       a   �  � � � �                             � � � �     c    ����     \�^�  � � � �       d   �  � � � �                             � � � �     f    ����     \�^�  X � h �       g   �  p � q �                             l � t �     i    ����                   ���  CWire�� 
 CCrossOver  ,4      m�  DL      m�  $      m�          � Y       k�  p!q      k�m�  4<        � 8�9     
 k�m�  \d      m�  4<      m�  ��      m�  ��      m�  ��      m�  ��      m�  |�        Xq       k�m�  \d        � `!a      k�m�  .,44      m�  .�4�      m�  .�4�      m�  .�4�      m�  .�4�      m�  .|4�      m�  .T4\      m�  .D4L      m�  .4$      m�  .4        0� 1       k�m�  ��      m�  � �� �      m�  .�4�        � �Q�      k�m�  ��      m�  � �� �      m�  .�4�        � �Q�      k�m�  ��      m�  � �� �      m�  � �� �      m�  .�4�      m�  � �� �      m�  � �� �        p �Q�      k�m�  ��      m�  � �� �      m�  .�4�        � �Q�      k�m�  |�      m�  � |� �      m�  � |� �      m�  .|4�      m�  � |� �      m�  � |� �        p �Q�      k�m�  � �� �      m�  � |� �        � H� a       k�m�  � �� �      m�  � �� �      m�  � �� �      m�  � �� �      m�  � |� �      m�  � D� L        � 0� 9      
 k�   �!1       k�   �!�       k�  ��!�      k�m�  � D� L      m�  .D4L      m�  � D� L      m�  � D� L      m�  DL        � HII      k�m�  ,4      m�  .,44        � 0�1     
 k�  �0�Q      
 k�  �(�)      k�m�  ����        ���)       k�  ����      k�m�  ����        ����      k�  ����      k�  ����       k�  �P�Q     
 k�  ����       k�  0 Q      k�m�  .T4\        XIY      k�m�  .4$      m�  $        �  I!      k�m�  � �� �      m�  � |� �      m�  � D� L      m�  � �         � � � �       k�m�  � �� �        � �� �       k�m�  � |� �      m�  � D� L        �  � �       k�m�  .4      m�  � �       m�        m�  � �       m�  � �         p I      k�m�  � �         � � � I       k�  p �q �       k�  ��     	 k�  ��      	 k�  ��     	 k�  � �Y       k�  �`��       k�  ����      k�  p q �       k�m�  � �         � � � !       k�  p � q        k�  0� 1�        k�  � 1�       k�  � � � �        k�  � � � �                     �                                      (  ! - ! # E # & } & ' r ' ( (  + � + , � , - - ! / � / 0 0 3 3 0 3 4 s 4 5 5 � 7 � 7 8 � 8 9 9 � ; � ; < � < = = � ? � ? @ � @ A A � C � C D � D E E # G � G H � H I I � K � K L � L M M � O � O P � P Q Q � S � S T � T U U � W � W X X  Z � Z [ [ � ` ` � c c � f f � i i � l � l � l � l � ` � u ' s w � 4 u ~ u t u � u � u � u � u � l r } v � &  �  �  �  �  �  �  �  �  �  � X � � x � � � � � ; � y � � � � � @ � z � � � � � � � � � � � ? � { � � � � � H � | � � � � � � � � � � � G � � � � � } � � � � � � � � � � � � � s , 5 � + 9 � � � � � � � � � � o � O � n � � � � � � � / � � � � A � � � = � � � 8 � Q K � 7  < � � u P � � � p � T � � � � � � � � [ � � � � � � � � � � � � � � � � q � � � � � S � � f � � � � C � � U � D M L � I � � � � � c � i � � W l � � Z � �             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 