��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  9�W    X1X4      �  9�[�    X2'X3'      �  9Y]g    X2+X3      �  9� [�     X1'X4'                    ��� 	 CLogicOut�� 	 CTerminal  �0�E       	        �            �D�T          ��    ��  \q      	        �            L\          ��    ��   ��      	       @            �$�          ��    ��  CNOR�  ����               �          �  ����               �          �  ���              @            ����           ��    ��  COR�  p(�)               �          �  p8�9               �          �  �0�1               �            �$�<           ��    ��  CAND�  0xEy               �          �  0�E�     	          �          �  \�q�               �            Dt\�     !      ��    ��  �`�a              @          �  �p�q                          �  �hi               �            �\�t     %      ��    ��  ��	               �          �  ��               �          �  �               �            ��     )      ��    ��  CXOR�  �0�1              @          �  �@�A              @          �  �8�9               �            �,�D     .      ��    ��  �h�i               �          �  �x�y               �          �  �pq               �            �d�|     2      ��    ��  � �!     	          �          �  �0�1     
         @          �  �(�)               �            ��4     6      ��    ��  ����               �          �  ����              @          �  ����               �            ����     :      ��    ��  (�=�              @          �  (�=�              @          �  T�i�              @            <�T�     >      ��    ��  (�=�               �          �  (�=�              @          �  T�i�               �            <�T�     B      ��    ,��  (@=A              @          �  (P=Q                          �  THiI     
         @            <<TT     F      ��    ��  ( =               �          �  (=               �          �  Ti	     	          �            <� T     J      ��    ��  CLogicIn�� 	 CLatchKey  0 � @ �      N   �  H � I �               @            D � L �     Q   ����     M�O�  ` � p �      R   �  x � y �               @            t � | �     T   ����     M�O�  � � � �       U   �  � � � �                             � � � �     W    ����     M�O�  � � � �      X   �  � � � �               @            � � � �     Z   ����     �� 	 CInverter�  ` � a �                @          �  ` � a �                �            T � l �     ]      ��    [��  � � � �                @          �  � � � �                �            � � � �     `      ��    [��  � � � �                            �  � � � �               @            � � � �     c      ��    [��  � 	�                @          �  � 	�                �            � � �     f      ��                  ���  CWire  q      i�  p�q      i�  ����      i�  ���1       i�  �p��       i�  p8q�       i�  pq)       i�  h�	     	 i�  �� �	      	 i��� 
 CCrossOver  � �       t�  � � � �       t�  � � � �       t�  � � � �       t�  � � � �       t�  v � | �       t�  ^ � d �       t�  F � L �         ( � ��      	 i�  ( � ) �      	 i�t�  � �       t�  �         � 	       i�t�  � � � �       t�  � �� �      t�  � �� �      t�  � �� �      t�  � L� T      t�  � <� D      t�  � � �         � � � �       i�t�  � � � �       t�  � �� �      t�  � L� T      t�  � <� D      t�  � � �         � � � �       i�t�  � � � �       t�  � <� D      t�  � � �         � � � Q       i�t�  � � � �       t�  � <� D      t�  � � �         � � � �       i�t�  v � | �       t�  v � |         x � y A       i�t�  ^ � d �         ` � a        i�t�  F � L �         H � I �       i�  ( �1�     	 i�  0h1y       i�  h1i      i�  � p�q      i�t�  � \� d      t�  � ,� 4      t�  � �� �      t�  � �� �        � P� q       i�t�  � \� d        x `�a      i�t�  � �� �      t�  v �| �      t�  � �� �        H �)�      i�t�  v ,| 4      t�  v �| �        x @y a       i�t�  � ,� 4      t�  v ,| 4      t�  � ,� 4        H 0�1      i�  � @�A      i�t�  v�|�        x�y	       i�  ��!      	 i�  x�	      i�t�  v�|�        h���      i�  h�y�      i�  h�i�       i�  ��9       i�  �8�9      i�t�  � ,� 4        � �� A       i�  H �I 1       i�  �x��       i�  ����      i�  �h�i      i�  �(�i       i�  ����       i�  ����       i�  h���      i�  �0�I      
 i�  hH�I     
 i�t�  � �� �        � �)�      i�t�  � � �       t�  � � �       t�  � � �       t�  � � �       t�  v � |       t�  �         `  )      i�t�  � �� �      t�  � �� �      t�  � �� �        � �)�      i�t�  � L� T      t�  � L� T        � P)Q      i�t�  � <� D      t�  � <� D      t�  � <� D      t�  � <� D        x @)A      i�  � �)�      i�  )      i�  H � a �       i�  ` � a �        i�  x � � �       i�  � � � �        i�  � � � �       i�  � � � �        i�  � � 	�       i�  � 	�                      �                                 4     n   l      p   o    m ! � ! " � " # # o % � % & � & ' ' � ) � ) * � * + + j . � . / � / 0 0 � 2 � 2 3 � 3 4 4 k 6 � 6 7 � 7 8 8 � : � : ; � ; < < � > � > ? � ? @ @ � B � B C � C D D � F � F G � G H H � J � J K � K L L q Q Q � T T � W W � Z Z � ] � ] ^ ^ � ` � ` a a � c � c d d � f � f g g ~ + p  n m  l  k   # j  L � s q s  s � s � s � s � s � s � s � } r s � ~ u ~ � g � � v � � � � � � � � � � � � Z � � w � � � � � � � � d � � x � � � � W � � y � � � � a � � z � � T � � { ^ � � | Q � } " � ! ' � � & � � � � � � � � � � � � � % � � � � � � � > � � � � � � � � � � � � � . � / � � � � r 6 � ) � � @ � � � D � * � 0 � � � � � � � 3 � < � � 2 8 � ; � � : � � 7 � H � � � � C � � � � � � � � � � � � � J � � � � � � � B � � � � � G � � � � � � � � � F � ? ~ K � � � ] � � � ` � � � c � � � f             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 