��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel   ! " /     X1      �  i ! z /     X2      �  � ! � /     X3      �  ! /     X4                  ��� 	 CInverter�� 	 CTerminal  �� ��               @          �  �� ��                �            �� ��            ��    ��  CAND�   � 5�                �          �   � 5�                �          �  L� a�                �            4� L�            ��    �� 	 CLogicOut�  �X�Y              @            �P�`          ��    ��  COR�  x�	              @          �  x�     
          �          �  ��              @            ��           ��    ��  x� ��               @          �  x� ��                �          �  �� ��               @            �� ��             ��    ��  (@=A               �          �  (P=Q                          �  THiI     
          �            <<TT     $      ��    ��  x@�A                          �  �@�A     	         @            �4�L     (      ��    ��  x �!              @          �  � �!               �            ��,     +      ��    ��  �(�)               �          �  �8�9     	         @          �  0!1               �            �$<     .      ��    ��  �� ��                           �  �� ��               @            �� ��      2      ��    ��  �� ��                           �  �� ��               @          �  � �                �            �� �      5      ��    ��  p %q               @          �  � %�               @          �  <x Qy               @            $l <�      9      ��    ��  CLogicIn�� 	 CLatchKey  �! �/      =   �  �, �A               @            �$ �,     @   ����     <�>�  ) (7       A   �  04 1I                             ,, 44     C    ����     <�>�  h) x7       D   �  �4 �I                             |, �4     F    ����     <�>�  �) �7      G   �  �4 �I               @            �, �4     I   ����     <�>�    A 0 O       J   �  8 L 9 a                             4 D < L     L    ����     <�>�  h A x O       M   �  � L � a                             | D � L     O    ����     <�>�  � A � O      P   �  � L � a               @            � D � L     R   ����     <�>�  � I  W       S   �  T 	i                             L T     U    ����     ��  0� E�                           �  \� q�               @            D� \�      W      ��    ��  0� E�                           �  \� q�               @            D� \�      Z      ��    ��  @hUi                          �  lh�i              @            T\lt     ]      ��    ��  @�U�              @          �  l���               �            T|l�     `      ��                ���  CWire�� 
 CCrossOver  � d� l        � hAi      c�  �� �       c�  �� ��        c�e�  ~� ��         `� ��       c�e�  ~� ��       e�  ~� ��       e�  ~l �t         �H ��        c�e�  ^� d�         `� a�        c�e�  ~� ��         `� ��       c�e�  ^� d�       e�  ~� ��         0� ��       c�e�  ~� ��         �� �       c�   � !�        c�  �� !�       c�  x� y�        c�  `� y�       c�   � !�        c�  � !�       c�  xyI      
 c�  �p �!       c�  �8�Y       c�  �8�9      c�  ��9       c�  x� y	       c�  x� ��       c�  �� ��        c�  hHyI     
 c�  xx y�        c�  Px yy       c�e�  �l �t         �H ��        c�  (P)Y       c�  XX)Y      c�e�  V<\D      e�  V\$        X YY       c�e�  V<\D        0@yA      c�e�  V\$      e�  .4$        � y!      c�  X �      c�  (0)A       c�   0)1      c�  �8�A      	 c�  �@�A     	 c�e�  .4$        0� 1A       c�  � �)       c�  � �!      c�e�  .l 4t         0H 1�        c�  �� ��       c�  �� ��       c�e�  ~l �t       e�  .l 4t       e�  �l �t         �p q       c�  �@ �q        c�  � 1�       c�e�  ~ � � �       e�  � � � �       e�  � �         8 � 1�       c�  8 ` 9 �        c�e�  � �         h 	�        c�  � �A�      c�e�  ~ � � �         � ` � i       c�e�  � d� l      e�  � � � �         � ` � �                   �                         q    y  |   x    {  �   �   ~    �   �   ! z ! " " � $ � $ % � % & & � ( � ( ) ) � + � + , , � . � . / � / 0 0 � 2 � 2 3 3 � 5 s 5 6 � 6 7 7 } 9 � 9 : g : ; ; � @ @ � C C � F F k I I � L L � O O � R R � U U � W � W X X   Z � Z [ [   ] d ] ^ ^   ` � ` a a   d � � ] � : g i i l o h k j k u k � F � o t i q q w o  s p s m � 5 v r k �  y  x ! {  z }  7 |  � � � �  � �  � �  � � " � & ~ �   ; � � � I h % � � � � � � � � � � � � ( � � � �  + � v � $ 0 � / � ) � � � � � � . , � � � C s 3 6 v 2 � n � � � �  9 @ � � Z � � � � � � � W L � � � U � � ` � � O d � f � � R �             �$s�        @     +        @            @    "V  (      �8                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 