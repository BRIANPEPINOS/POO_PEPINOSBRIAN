��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  �%'    
X1X2'X3'X4      �  ���    X1'X4'+(X2xorX3)      �  Q� ��     X1XORX4      �  !� C�     X2'X3'      �  )�G�    X2X3      �  )AKO    X1'X4'                    ��� 	 CLogicOut�� 	 CTerminal  `�u�     % 	       @            t���          ��    ��  COR�   �5�               �          �   �5�     #         @          �  L�a�     %         @            4�L�           ��    �� 	 CInverter�  h(})               �          �  �(�)     $         @            |�4           ��    ��  CAND�  � �     "         @          �  ��     $         @          �  �		     #         @            ���           ��    ��  h }               �          �  � �     "         @            |��     "      ��    ��  �� ��                @          �  �� ��                �            |� ��     %      ��    ��  H� I�       !         @          �  H� I�                �            <� T�     (      ��    ��  � �                @          �  � �                �            � $�     +      ��    ��  �� ��                             �  �� ��               @            �� ��     .      ��    ��  CLogicIn�� 	 CLatchKey  Pa `o      1   �  hl i�               @            dd ll     4   ����     0�2�  a (o      5   �  0l 1�      !         @            ,d 4l     7   ����     0�2�  �a �o      8   �  �l ��               @            �d �l     :   ����     0�2�  �a �o       ;   �  �l ��                              �d �l     =    ����     ��  �� ��                            �  �� ��      !         @          �  �� ��                �            �� ��      ?      ��    ��  ��              @          �  � �!              @          �  ��              @            ��$     C      ��    ��  �H�I              @          �  �X�Y               �          �  �P�Q               �            �D�\     G      ��    ��  �x�y               �          �  ����               �          �  ����               �            �t��     K      ��    ��  �`a               �          �  �pq               �          �  h1i               �            \t     O      ��    ��   � �                �          �   	              @          �  , A              @            � ,     S      ��    ��  H(])              @          �  H8]9               �          �  t0�1              @            \$t<     W      ��    ��  ��1      	       @            ��    [     ��    ��  ����               �          �  ����              @          �  ����               �            ����     ]      ��    ��  CXOR�   �5�                          �   �5�              @          �  L�a�              @            4�L�     b      ��    ��   -              @          �  -               �          �  DY	     	          �            ,� D     f      ��    ��  �-�                          �  �-�              @          �  D�Y�               �            ,|D�     j      ��    ��  X-Y              @          �  h-i               �          �  D`Ya               �            ,TDl     n      ��    ��  (4)I      	        �             $04    r      ��    ��  �@�A               �          �  �P�Q               �          �  H)I               �            �<T     t      ��    ��  `hui               �          �  `xuy               �          �  �p�q               �            td�|     x      ��    ��  �� ��      	          �          �  ��	               �          �  � �               �            �� �     |      ��    ��  `0u1     
         @          �  �0�1               �            t$�<     �      ��    `��  (-)                          �  8-9              @          �  D0Y1     
         @            ,$D<     �      ��    ��  � � � �                @          �  � � � �                �            � � � �     �      ��    ��  � � � �                @          �  � � � �                �            � � � �     �      ��    ��  � � � �                            �  � � � �               @            t � � �     �      ��    ��  H � I �                            �  H � I �               @            < � T �     �      ��    0�2�  � � � �      �   �  � � � �               @            � � � �     �   ����     0�2�  � � � �      �   �  � � � �               @            � � � �     �   ����     0�2�  H � X �       �   �  ` � a �                             \ � d �     �    ����     0�2�   � ( �       �   �  0 � 1 �                             , � 4 �     �    ����                   ���  CWire�� 
 CCrossOver  � �� �        ` �!�      ��  � �!�      ��  X�Y�       ����  ����        ����       ����  � �� �        � �� �       ��   �!	      # ��  !	     # ��   �!�       ��  ��!�      ��  ��     $ ��  ��)      $ ��  P(i)      ��  P�Q)       ����  n�t�        P���      ����  n�t�      ��  n�t�        p�q�       ��  ����      ����  ����      ��  n�t�        `���      ����  �L�T        �H��       ��  � �     " ��  h�i       ��  h�q�      ��  X�q�      ��  �� ��        ��  h� ��       ��  H� I�       ! ��  � �        ��  �� ��         ��  �� ��        ��  �� ��         ��  0� I�      ! ��  �� �       ����  fl      ��  f� l�       ��  f� l�         h� i!       ����  �� ��         �� �       ����  �� ��         �� �I       ����  .� 4�         0� 1�       ! ����  DL      ��        ��  � �         � Y       ����  FTL\      ��  FDLL      ��  FL      ��  F� L�       ��  F� L�         H� Iy       ����  �� ��       ��  F� L�       ��  � �       ��  �� ��       ��  f� l�       ��  �� ��       ��  .� 4�         �� ��        ����  �� ��       ��  F� L�       ��  f� l�         0� ��      ! ����  ��      ��  FL      ��        ��  fl        ��      ����  ��$        h �!      ����  �D�L      ��  FDLL      ��  DL        �H�I      ����  �T�\      ��  FTL\        X�Y      ����  �t�|        Hx�y      ����  �t�|      ��  �T�\      ��  �D�L      ��  ��$      ��  ��      ��  �� ��       ��  �� ��         �� ��       ��  ����      ��  �P�a       ��  �p��       ��  �� �       ��   � �        ��  �      ��          ��  @ A)       ��  @(I)      ��  081i       ��  08I9      ��  �P�q       ����  �L�T        �P�Q      ��  XH�I      ��  XHYa       ��  ����       ��  ` �a �       ��  �� ��      	 ��  �� �	      	 ��  X�	     	 ����  � �         �       ����  � � �         � � �        ����  � �       ��  � � �       ��  � $� ,      ��  � 4� <      ��  � T� \        � � � i       ����  � � �       ��  � � �       ��  � � �         �        ��  � � �        ����  � � �       ��  � $� ,        � � � 9       ����  ^ $d ,      ��  � $� ,      ��  F $L ,      ��  � $� ,        0 ()      ����  ^ Td \      ��  ^ $d ,        ` � a �       ��  Xxay      ��  XxY�       ��  Xhai      ��  X`Yi       ��  � ��      ����  � |� �      ��  � T� \        � 8� �       ����  � |� �        ` ��      ����  � T� \      ��  ^ Td \      ��  � T� \        H XY      ��  � hi      ����  � 4� <        � 89      ����  F $L ,        H � I Y       ��  �@�A      ��  � �A       ��  ��1       ��  X0a1     
 ��  0 � 1 )       ��  � � � �        ��  � � � �       ��  � � � �        ��  � � � �       ��  � � � �        ��  ` � � �       ��  H � I �        ��  0 � I �                     �                                �   �      �    �  �   �      � " � " # # � % � % & & � ( � ( ) ) � + � + , , � . � . / / � 4 4 � 7 7 � : : � = = � ? � ? @ � @ A A C � C D � D E E G � G H � H I I K � K L L M M O O P P Q Q 
S S T T U U W 	W X X Y Y [ [ [ Y ] � ] ^ ^ _ _ � b � b c � c d d � f  f g g h h j 8j k 4k l l 1n :n o >o p p r r v t Ct u u v v r x 2x y 0y z z | | } E} ~ ~ D� F� � � E� (� � ?� � � F� H� � � � J� � � � L� � � $� N� � � A� � I� � K� � M� � O� � b � c l � � � � � � � 4�  �   � �  _ � �  �  �  � � � � � � � � � � � � � ] � � � � d � � #  � " � � � � � % � � � ( � + � . � � = � � � � � � � � � � � 4 � � � : � � � / � � � 7 � � � � � � � , � � � � � � � � � � � ) � �  � � � � � � � � � � � � � ? � � � � � � � @ � � � � � � � � � C � � � D � � � � � � � G � � � � � H � � � K � � � � � � � � � � � � � � & � L I O P M A S E T U 	W Q 
X z � u � 3^ � -� | h g !� "*@=� >   &$f �  %#%,� 5(/((B('G� -<-)� 81y 0� 3x p 25k 595;?� 86j :7:.:An o ?%� A+� :Dt ~ C} � � � � (I� � HK� %JM� -LO� GN &           �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 