��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  ��8     F(A,B,C)=A'B'C'+A'BC'+AB'C'+ABC'      �  	�O�    (A'BC')+(ABC')      �  ��C�    (A'B'C')+(AB'C')      �  ����    ABC'      �  �A�O    A'BC'      �  I!]/    BC'      �  I�f�    AB'C'      �  Q�p�    A'B'C'      �  aQn_    C'      �  �I�W    B'C'      �  � Q� _    A'      �  Q&_    B'      �  )� 4�     C      �  � � � �     B      �  I � T �     A      �  i � �      F(A,B,C)=A'B'C'+A'BC'+AB'C'+ABC'                    ��� 	 CLogicOut�� 	 CTerminal  �(�)      	        �            � �0           ��    ��  COR�  P e!               �          �  P0e1               �          �  |(�)               �            d|4           ��    ��  ����               �          �  ����               �          �  �!�               �            ���     #      ��    ��  ����               �          �  ����     	          �          �  ��               �            ���     '      ��    ��  CAND�  p���     
          �          �  p���              @          �  ����               �            ����     ,      ��    *��  �`�a     
          �          �  �p�q               �          �  �h�i               �            �\�t     0      ��    *��  (�=�               �          �  (=	              @          �  T i     	          �            <�T     4      ��    *��  (8=9               �          �  (H=I              @          �  T@iA     
          �            <4TL     8      ��    *��  0�E�               �          �  0�E�               �          �  \�q�               �            D�\�     <      ��    *��  �p�q               �          �  ����               �          �  �xy               �            �l��     @      ��    �� 	 CInverter�  pq               @          �  p4qI               �            d|4    E      ��    C��  	               @          �  4	I               �            � 4    H      ��    C��  � �                @          �  � 4� I               �            � � 4    K      ��    ��  CLogicIn�� 	 CLatchKey  ` � p �      N   �  x � y �               @            t � | �     Q   ����     M�O�  � � � �      R   �  � � � �               @            � � � �     T   ����     M�O�  (� 8�      U   �  @� A�               @            <� D�     W   ����                   ���  CWire  P0Q�       Y�   �Q�      Y�  P�Q!       Y�  �Q�      Y�  ����       Y�  ����      Y�  �h��       Y�  �h�i      Y�  ���      	 Y�  h �     	 Y�  ����       Y�  p���      Y��� 
 CCrossOver  � �       g�  � �       g�  nt        x )	      Y�  x y �       Y�  x �q�      Y�g�  fllt        h@i�      
 Y�g�  fllt        � p�q      Y�  h�q�     
 Y�  h@�A     
 Y�g�  � �� �      g�  n�t�      g�  ���        � �1�      Y�g�  � �         � �� q       Y�g�  � �� �      g�  � �         � � � I       Y�  � H)I      Y�  �@�a      
 Y�  � � � 	       Y�  H	�       Y�  p8)9      Y�  pp�q      Y�g�  n|t�      g�  n�t�      g�  nt        ppq9       Y�g�  n|t�        ���      Y�  x � y 	       Y�g�  ���         x�       Y�   �)�      Y�  � H� �       Y�   x1y      Y�  0x1�       Y�  pHqq       Y�  p� q	       Y�  @� q�       Y�  � 		       Y�  � � 	�       Y�  x � � �                     �                             !   \    Z   ! !  # ` # $ ^ $ % % [ ' d ' ( b ( ) ) ] , q , - l - . . _ 0 } 0 1 o 1 2 2 a 4 � 4 5 f 5 6 6 c 8 � 8 9 | 9 : : r < � < = s = > > e @ � @ A � A B B � E � E F F � H � H I I  K ~ K L L � Q Q � T T � W W �   [ % Z ]  ) \ $ _ . ^ a # 2 ` ( c 6 b e ' > d f x f { f � � 5 f l k - m p : q o n w 1 m , m } s z s � s � � = w h s o y t y i T | y 9 r 0 � K I � � 8 � @ � � � u � j � � � �  A Q k � v B � � 4 L w � � � < F � � E W � � H y � � ~             �$s�        @     +        @            @    "V  (      �8                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 