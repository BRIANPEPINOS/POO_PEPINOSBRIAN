��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  ��    X2X3      �  �)(7    X1X3'X4'      �  ��(�    X1'X2'X4      �  I�y�    EMPATA      �  ����    GANA B      �  �� ��     GANA A      �  �0�    X1'X2'X3      �  I0W    X2X3'X4'      �  ����    X1'X2'      �  ����    X3'X4'      �  �	�    X1X4                    ��� 	 CLogicOut�� 	 CTerminal  �h�}       	        �            �|��          ��    ��  ��1      	        �            ��          ��    ��  8�M�      	       @            L�\�          ��    ��  CNOR�  ���               �          �  ���               �          �  $�9�              @            �$�           ��    ��  COR�  �`�a               �          �  �p�q               �          �  �h�i               �            �\�t     #      ��    !��  @ U!               �          �  @0U1               �          �  l(�)               �            Tl4     '      ��    ��  CAND�  �xy              @          �  ���                          �  �1�               �            t�     ,      ��    *��  �@A               �          �  �PQ                          �  H1I               �            <T     0      ��    *��  � �               �          �  ��              @          �  )	               �            ��     4      ��    !��  �(�)     	          �          �  �8�9               �          �  �0�1               �            �$�<     8      ��    !��  @�U�               �          �  @�U�               �          �  l���               �            T|l�     <      ��    *��  ���                          �  ���               �          �  �1�               �            ��     @      ��    *��  �`a              @          �  �pq               �          �  h1i               �            \t     D      ��    *��  ����              @          �  ����               �          �  ����               �            ����     H      ��    *��  �h�i              @          �  �x�y               �          �  �p�q               �            �d�|     L      ��    *��  �(�)                          �  �8�9              @          �  �0�1     	          �            �$�<     P      ��    �� 	 CInverter�  X� Y�                @          �  X� Y               �            L� d�     U      ��    S��  � �                            �  �               @            � $�     X      ��    S��  � � � �                @          �  � � �                �            � � � �     [      ��    S��  � � � �                            �  � � �               @            � � � �     ^      ��    ��  CLogicIn�� 	 CLatchKey   � 0�      a   �  8� 9�               @            4� <�     d   ����     `�b�  � � � �       e   �   � �                             � � �     g    ����     `�b�  � � � �      h   �  � � � �               @            � � � �     j   ����     `�b�  � � � �       k   �  � � � �                             � � � �     m    ����                   ���  CWire  �0�1      o�  �0��       o�  ���i       o�  �h�i      o�  �(�a       o�  �(�)      o�  �p��       o�  0���      o�  @0AI       o�  0HAI      o�  @A!       o�  (A	      o�   ���      o��� 
 CCrossOver  � t|      ~�  � LT      ~�  � ��      ~�  � ��         ��       o�~�  � t|        � x�y      o�~�  � LT      ~�  � L� T        � P�Q      o�~�  � ��      ~�  6�<�        � ���      o�~�  � L� T      ~�  � �� �        � X� y       o�~�  � ��      ~�  � �� �      ~�  6�<�      ~�  � �� �        � ���      o�  � (� Q       o�  �@�A      o�~�  ��      ~�  ���      ~�  ����      ~�  ����        �p�A       o�  �p�q      o�~�  ��        8�      o�~�  ���        � �      o�~�  ����        ����      o�~�  ����      ~�  6�<�        ���      o�  �p�q      o�~�  6�<�      ~�  6�<�      ~�  6�<�      ~�  6d<l      ~�  6T<\        889       o�~�  6d<l      ~�  Vd\l        h�i      o�~�  6T<\      ~�  � T\      ~�  VT\\      ~�  T\      ~�  � T� \        � X�Y      o�  ���       o�  ����      o�  �8��       o�  �(�1      	 o�  �0�1     	 o�  @�A�       o�  0�A�      o�  @hA�       o�  0hAi      o�  ����       o�  �	�       o�   �	�      o�~�  � T\      ~�  � $,         � �       o�~�  � $,      ~�  � $� ,      ~�  � $� ,      ~�  � $� ,      ~�  V$\,      ~�  $,      ~�  6$<,        � (�)      o�  �X�a       o�~�  � $� ,        � � � Y       o�~�  VT\\      ~�  Vd\l      ~�  V4\<      ~�  V$\,        XYy       o�~�  T\      ~�  $,        i       o�~�  � T� \      ~�  � �� �      ~�  � $� ,        � � �       o�~�  � $� ,        � � �       o�  Xx�y      o�~�  V4\<        88�9      o�  � � � )       o�~�  6$<,        8� 99       o�  X� Y�        o�  8� Y�       o�  � �        o�   � �       o�  � � � �        o�  � � � �       o�  � � � �        o�  � � � �                     �                             %    :      q   r       # t # $ v $ % % s ' z ' ( x ( ) ) u , � , - | - . . w 0 � 0 1 � 1 2 2 y 4 � 4 5 � 5 6 6 { 8 � 8 9 � 9 : : p < � < = � = > > � @ � @ A � A B B � D � D E � E F F � H � H I � I J J � L � L M � M N N � P � P Q � Q R R � U � U V V � X � X Y Y � [ � [ \ \ � ^ � ^ _ _ � d d � g g � j j � m m �  q p   s  r u # ) t $ w . v ( y 2 x { ' 6 z } - } � } � } � } � � | �  � , � � � � � 1 � � � � � I � � � � � � � � � � � � � � � H � � � 0 � � � � � � � � � � N � � � � 5 � � � 4 � � � A � � � � � � � E � � � � � � � � � � � � � � � � � L � � � � � � � � � � � � J � > � 9 � 8 � R � = � B � � < F � � @ � � � � � � � � g } � � � � � � � � � � � � � � � P � D � � j � � � � � � � � � V � � � � � Y � � � � � � � \ � � � _ � � M � � � Q m � � � � � � U d � � X � � � [ � � � ^ � �             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 