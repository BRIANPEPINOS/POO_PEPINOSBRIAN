��  CCircuit��  CSerializeHack           ��  CPart    �   �     ��� 	 CLogicOut�� 	 CTerminal  PQ              @            H�X         ��    ��  CAND
�  Ppeq                          
�  P�e�               �          
�  |x�y               �            dl|�           ��    �
�  ����               �          
�  ����               �          
�  ����               �            ����           ��    �
�  �@�A              @          
�  �P�Q              @          
�  �H�I              @            �<�T           ��    �
�  Pe              @          
�  P e!              @          
�  |�              @            d|$           ��    �
�  P�e�                          
�  P�e�              @          
�  |���               �            d�|�           ��    ��  CLogicIn�� 	 CLatchKey   AO      "   
�  La                            DL    %    ����     !�#�  PA`O      &   
�  hLia                            dDlL    (    ����     !�#�  �A�O     )   
�  �L�a              @            �D�L    +   ����     !�#�  �AO     ,   
�  La              @            DL    .   ����     �� 	 CInverter
�  0p1�                           
�  0�1�              @            $�<�    1      ��    /�
�  �x��                           
�  ����              @            t���    4      ��    /�
�  �x��               @          
�  ����               �            ����    7      ��    /�
�  0x1�               @          
�  0�1�               �            $�<�    :      ��    ��  COR
�  � �               �          
�  ��              @          
�  	              @            ��     >      ��    <�
�  `a              @          
�  pq               �          
�  4hIi              @            \4t     B      ��    �
�  h }              @          
�  h}                          
�  ��	     
          �            |� �     F      ��    �
�  @� U�       	        �            T� d�      J      ��    <�
�   � �                �          
�   � �                �          
�  ,� A�                �            � ,�      L      ��    �
�  � �!     
          �          
�  �0�1               �          
�  �(�)               �            ��4     P      ��    �
�  �� ��                �          
�  �� ��               @          
�  �� ��                �            �� ��      T      ��    ��  CXOR
�  `� u�                           
�  `� u�               @          
�  �� ��               @            t� ��      Y      ��    �
�  h@}A              @          
�  hP}Q     	          �          
�  �H�I               �            |<�T     ]      ��    �
�  `� u�               @          
�  `� u�                �          
�  �� ��                �            t� ��      a      ��    /�
�  8@ 9U                @          
�  8l 9�      	          �            ,T Dl     e      ��    /�
�  � @ � U                @          
�  � l � �                �            � T � l     h      ��    /�
�  � @ � U                            
�  � l � �               @            | T � l     k      ��    /�
�  8 8 9 M                            
�  8 d 9 y               @            , L D d     n      ��    !�#�   	       p   
�   )               @                  r   ����     !�#�  � 	 �       s   
�  �  � )               @            �  �      u   ����     !�#�  X 	 h        v   
�  p  q )                             l  t      x    ����     !�#�   	         y   
�     ! )                               $      {    ����         �   �     ���  CWire  HQ      }�  HIi       }�  ��A       }��� 
 CCrossOver  ~�      ��  ~���        ���!       }�  0�1       }�  `q       }�  �x��       }�  0���      }���  .|4�      ��  .l4t      ��  .L4T      ��  .4$      ��  .4      ��  .�4�      ��  .�4�        0�1�       }���  .|4�        ��Q�      }���  .l4t      ��  �l�t        pQq      }���  .L4T        P�Q      }���  .4      ��  ��      ��        ��  ~�        0Q      }���  .�4�      ��  ����      ��  ��        ��Q�      }���  .�4�      ��  ����      ��  ��      ��  ~���      ��  ����        h�Q�      }���  .4$      ��  ��$      ��  $        � Q!      }���  $      ��        ��  ��      ��  ��        `Q       }���  ����        �`��       }�  h`i�       }�  `1a      }�  0`1q       }�  h`�a      }�  �`�y       }�  `1a      }�  0`1y       }�  �`�y       }�  �`�a      }�  ��      }�  ����      }�  ���       }�  ��I       }�  I       }�   HI      }�   Ha       }�   `	a      }�  ��	�      }�  p	�       }���  �l�t      ��  ��$      ��  ��      ��  ����      ��  ����        ����       }�  � �!     
 }�  ��!      
 }���  6<      ��  � �         p i      }���  n � t       ��  n � t �         p ( q        }���  6<      ��  6� <      ��  6<<D      ��  6� <�       ��  6� <�       ��  6� <�       ��  6� <�         8� 9Q      	 }���  � �       ��  � � �       ��  � � � �       ��  � � � �         � ( � A       }���  n � t       ��  6� <      ��  � � �         8  i      }���  n � t �       ��  6 � < �       ��  6� <�       ��  � � � �       ��  � �           � a�       }���  6 � < �         8 x 9        }�  �� �       }�  �� �)       }�  �0�I       }�  �H�I      }�  �� �       }�  �� ��        }�  �� ��        }�  �� ��       }�  �� ��        }�  �� ��       }�  8PiQ     	 }���  6<<D        � @iA      }���  6� <�         � a�       }���  6� <�       ��  � �         � � a�       }���  6� <�       ��  � � � �       ��  � �       ��  � � � �         � � a�       }�  � ( � )       }���  � �       ��  � �       ��  � �         ( �        }�    ( ! �        }���  � � � �         � � � �        }�  � � � �        }�  � ( � A        }�  ( 9)       }�  � ( � A        }�  p ( � )       }�  8 ( 9 9        }�    ( 9 )       }�  8( 9A            �   �     �    �   �         �   �       ~  �   �    �  �   �    �  �   �    �  �   �    �  �   �      � % % � ( ( � + + � . . � 1 � 1 2 2 � 4 � 4 5 5 � 7 � 7 8 8 � : � : ; ; � > � > ? � ? @ @ � B � B C � C D D  F � F G � G H H � J N J L � L M � M N N J P � P Q � Q R R � T � T U � U V V � Y � Y Z � Z [ [ � ] � ] ^ � ^ _ _ � a � a b � b c c � e e f f � h h i i 	k k l l n n o o � r r u u x x { {   ~ D   � � � � 5 � 2 � % �   �  � � � � � � � � � � � � � � ; � � � �  � � � � �  � � �  � � � � � � � � �  � � � � � � �  � � � � � � � � � � �  � � � � � � �  � � � � � � � � . � � � + � ( � � � � 1 � � � 7 � � � : � 4 � � � ?   � � > �  @ � � � � � � B  � C � � � � � � � � � � � 8 � � P H � � � � � � G � � � � x � � � � � � � � � � � � � � � f � � � � � � � �  u � � � � � � � � F � � � � � � � � � Y � � o � � M � R Q � _ � � L V � U � [ � � T c � � ^ � � � ] � � Z � � � 	b � � � � � � 
a � � � r � { � 	i � l � k h � n e             �$s�        @     +        @            @    "V  (      ��                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 